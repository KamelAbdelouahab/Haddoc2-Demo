library ieee;
	use	ieee.std_logic_1164.all;
	use	ieee.numeric_std.all;

entity cnn_slave is
end cnn_slave;

architecture rtl of cnn_slave is
begin
end rtl;
